-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "11/12/2023 18:53:46"
                                                            
-- Vhdl Test Bench template for design  :  counting
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;                                               
USE ieee.std_logic_1164.all;                                

ENTITY counting_vhd_tst IS
END counting_vhd_tst;
ARCHITECTURE counting_arch OF counting_vhd_tst IS
-- constants                                                 
-- signals                                                   
SIGNAL clk_50M : STD_LOGIC;
SIGNAL continu : STD_LOGIC;
SIGNAL data_anemometre : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL data_valid : STD_LOGIC;
SIGNAL freq_in : STD_LOGIC;
SIGNAL reset : STD_LOGIC;
SIGNAL start_stop : STD_LOGIC;
COMPONENT counting
	PORT (
	clk_50M : IN STD_LOGIC;
	continu : IN STD_LOGIC;
	data_anemometre : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data_valid : OUT STD_LOGIC;
	freq_in : IN STD_LOGIC;
	reset : IN STD_LOGIC;
	start_stop : IN STD_LOGIC
	);
END COMPONENT;
BEGIN
	i1 : counting
	PORT MAP (
-- list connections between master ports and signals
	clk_50M => clk_50M,
	continu => continu,
	data_anemometre => data_anemometre,
	data_valid => data_valid,
	freq_in => freq_in,
	reset => reset,
	start_stop => start_stop
	);
clk_stimulus : process
begin
   wait for 10 ns;
		clk_50M <= not clk_50M;
end process clk_stimulus;

in_freq_anemometre_stimulus : process
begin

	wait for 500 ms;
	freq_in <= not freq_in;
end process in_freq_anemometre_stimulus;                                          
END counting_arch;
