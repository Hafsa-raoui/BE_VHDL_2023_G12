-------------------------------- LIBRARIES -----------------------------
library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-------------------------------- ENTITY ---------------------------
entity pwm is
	port(
		-- entree
		clk			: in std_logic;
		freq 		: in std_logic_vector (7 downto 0);
		duty		: in std_logic_vector(7 downto 0);
		reset		: in std_logic;
		-- sortie
		pwm_out		: out std_logic
		);
end pwm ;

--------------------------------- ARCHITRECTURE ------------------------
architecture arch of pwm is
signal count : std_logic_vector (7 downto 0);
begin
process(clk)
variable cpt : integer range 0 to 50000001; -- On a une horloge de fr�quence 50MHz donc 50000000 front montant pour une p�riode

begin
if reset='1' then pwm_out <='0'; -- Reset actif

else if (clk'event and clk='1') then
	cpt := cpt + 1 ;
	if  cpt <= duty then
		pwm_out <= '1';
	else if(cpt>= duty and cpt < freq-1) then 
		pwm_out <= '0';
	end if;
	if cpt = freq then
		cpt := 0;
	end if;
	
	end if;
	end if;
	
end if;

end process;
	
end arch;































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































